module tx(
    // Inputs
    input s_tick, clk, reset, tx_start,
    input [7:0] din,
    // Outputs
    output reg tx,
    output reg tx_done_tick
);


endmodule